`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:58:12 03/26/2017
// Design Name:   encoder8_3_2
// Module Name:   C:/Users/zhenyu/Documents/ise/system/encoder8_3/encoder8_3_2/encoder_8_3_2test.v
// Project Name:  encoder8_3_2
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: encoder8_3_2
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module encoder_8_3_2test;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	encoder8_3_2 uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

